`timescale 1ns/1ps

// Integration step 1: CSR + Command Engine
// - Verifies CMD_TRIGGER path, trigger clear, and CE latching
// - Checks PSLVERR behavior when busy, and XIP exclusivity
module int_csr_ce_tb;
  // Clock/reset
  reg clk; reg resetn;

  // APB
  reg        psel; reg penable; reg pwrite; reg [11:0] paddr; reg [31:0] pwdata; reg [3:0] pstrb;
  wire [31:0] prdata; wire pready; wire pslverr;

  // CSR <-> CE wires
  wire enable_w, xip_en_w, quad_en_w, cpol_w, cpha_w, lsb_first_w, cmd_start_w, dma_en_w, mode_en_w;
  wire hold_en_w, wp_en_w; wire [2:0] clk_div_w; wire cs_auto_w; wire [1:0] cs_level_w, cs_delay_w;
  wire [1:0] cmd_lanes_w, addr_lanes_w, data_lanes_w, addr_bytes_w; wire [3:0] dummy_cycles_w;
  wire is_write_w; wire [7:0] opcode_w, mode_bits_w; wire [31:0] cmd_addr_w, cmd_len_w; wire [7:0] extra_dummy_w;
  wire [3:0] burst_size_w; wire dma_dir_w; wire incr_addr_w; wire [31:0] dma_addr_w, dma_len_w;
  wire [31:0] fifo_tx_data_csr_w; wire fifo_tx_we_csr_w; wire [31:0] fifo_rx_rd_data_w; wire fifo_rx_re_csr_w;
  wire [4:0] int_en_w;
  wire cmd_trigger_clr_w;

  // CE wires
  wire ce_start_w, ce_busy_w, ce_cmd_done_set_w;

  // ID/status taps
  wire [31:0] csr_status_w;

  // CSR
  csr u_csr (
    .pclk(clk), .presetn(resetn),
    .psel(psel), .penable(penable), .pwrite(pwrite), .paddr(paddr), .pwdata(pwdata), .pstrb(pstrb),
    .prdata(prdata), .pready(pready), .pslverr(pslverr),
    .enable_o(enable_w), .xip_en_o(xip_en_w), .quad_en_o(quad_en_w), .cpol_o(cpol_w), .cpha_o(cpha_w), .lsb_first_o(lsb_first_w),
    .cmd_start_o(cmd_start_w), .dma_en_o(dma_en_w), .mode_en_o(mode_en_w), .hold_en_o(hold_en_w), .wp_en_o(wp_en_w),
    .cmd_trigger_clr_i(cmd_trigger_clr_w),
    .clk_div_o(clk_div_w), .cs_auto_o(cs_auto_w), .cs_level_o(cs_level_w), .cs_delay_o(cs_delay_w),
    .xip_addr_bytes_o(), .xip_data_lanes_o(), .xip_dummy_cycles_o(), .xip_cont_read_o(), .xip_mode_en_o(), .xip_write_en_o(),
    .xip_read_op_o(), .xip_mode_bits_o(), .xip_write_op_o(),
    .cmd_lanes_o(cmd_lanes_w), .addr_lanes_o(addr_lanes_w), .data_lanes_o(data_lanes_w), .addr_bytes_o(addr_bytes_w),
    .mode_en_cfg_o(), .dummy_cycles_o(dummy_cycles_w), .is_write_o(is_write_w), .opcode_o(opcode_w), .mode_bits_o(mode_bits_w),
    .cmd_addr_o(cmd_addr_w), .cmd_len_o(cmd_len_w), .extra_dummy_o(extra_dummy_w),
    .burst_size_o(burst_size_w), .dma_dir_o(dma_dir_w), .incr_addr_o(incr_addr_w), .dma_addr_o(dma_addr_w), .dma_len_o(dma_len_w),
    .fifo_tx_data_o(fifo_tx_data_csr_w), .fifo_tx_we_o(fifo_tx_we_csr_w), .fifo_rx_data_i(32'h0), .fifo_rx_re_o(fifo_rx_re_csr_w),
    .int_en_o(int_en_w),
    .cmd_done_set_i(ce_cmd_done_set_w), .dma_done_set_i(1'b0), .err_set_i(1'b0), .fifo_tx_empty_set_i(1'b0), .fifo_rx_full_set_i(1'b0),
    .busy_i(ce_busy_w), .xip_active_i(1'b0), .cmd_done_i(1'b0), .dma_done_i(1'b0),
    .tx_level_i(4'h0), .rx_level_i(4'h0), .tx_empty_i(1'b1), .rx_full_i(1'b0),
    .timeout_i(1'b0), .overrun_i(1'b0), .underrun_i(1'b0), .axi_err_i(1'b0), .irq()
  );

  // CE
  reg ce_done_i;
  cmd_engine #(.ADDR_WIDTH(32)) u_ce (
    .clk(clk), .resetn(resetn),
    .cmd_start_i(cmd_start_w), .cmd_trigger_clr_o(cmd_trigger_clr_w), .cmd_done_set_o(ce_cmd_done_set_w), .busy_o(ce_busy_w),
    .cmd_lanes_i(cmd_lanes_w), .addr_lanes_i(addr_lanes_w), .data_lanes_i(data_lanes_w), .addr_bytes_i(addr_bytes_w),
    .mode_en_i(mode_en_w), .dummy_cycles_i(dummy_cycles_w), .extra_dummy_i(extra_dummy_w), .is_write_i(is_write_w),
    .opcode_i(opcode_w), .mode_bits_i(mode_bits_w), .cmd_addr_i(cmd_addr_w), .cmd_len_i(cmd_len_w),
    .quad_en_i(quad_en_w), .cs_auto_i(cs_auto_w), .xip_cont_read_i(1'b0), .clk_div_i(clk_div_w), .cpol_i(cpol_w), .cpha_i(cpha_w),
    .start_o(ce_start_w), .done_i(ce_done_i),
    .cmd_lanes_o(), .addr_lanes_o(), .data_lanes_o(), .addr_bytes_o(), .mode_en_o(), .dummy_cycles_o(), .dir_o(),
    .quad_en_o(), .cs_auto_o(), .xip_cont_read_o(), .opcode_o(), .mode_bits_o(), .addr_o(), .len_o(), .clk_div_o(), .cpol_o(), .cpha_o()
  );

  // Clocking
  initial clk=0; always #5 clk=~clk; initial resetn=0;

  // APB helpers
  task apb_write(input [11:0] addr, input [31:0] data);
  begin @(posedge clk); psel<=1;penable<=0;pwrite<=1;paddr<=addr;pwdata<=data;pstrb<=4'hF; @(posedge clk); penable<=1; @(posedge clk);
        psel<=0;penable<=0;pwrite<=0;paddr<=0;pwdata<=0;pstrb<=0; end endtask
  task apb_read(input [11:0] addr, output [31:0] data);
  begin @(posedge clk); psel<=1;penable<=0;pwrite<=0;paddr<=addr; @(posedge clk); penable<=1; @(posedge clk); data=prdata; psel<=0; penable<=0; paddr<=0; end endtask

  // CSR addrs
  localparam CTRL=12'h004, CMD_CFG=12'h024, CMD_OP=12'h028, CMD_ADDR=12'h02C, CMD_LEN=12'h030;

  // Test
  initial begin
    psel=0;penable=0;pwrite=0;paddr=0;pwdata=0;pstrb=0; ce_done_i=0; repeat(5) @(posedge clk); resetn=1;

    // Enable controller and set Mode0
    apb_write(CTRL, 32'h0000_0001);
    // Configure 0x03 read 4B @ 0, 3B addr
    apb_write(CMD_CFG, 32'h0000_0040);
    apb_write(CMD_OP,  32'h0000_0003);
    apb_write(CMD_ADDR,32'h0000_0000);
    apb_write(CMD_LEN, 32'h0000_0004);
    // Trigger
    apb_write(CTRL, 32'h0000_0101);
    // CE should assert start then we complete it
    repeat(4) @(posedge clk); ce_done_i<=1; @(posedge clk); ce_done_i<=0;
    repeat(4) @(posedge clk);
    $display("CSR+CE integration test passed");
    $finish;
  end

  // Global timeout to prevent stalls
  initial begin
    #1_000_000; // 1 ms cutoff
    $display("[int_csr_ce_tb] Global timeout reached — finishing.");
    $finish;
  end
endmodule
