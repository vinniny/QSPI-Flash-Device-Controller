`timescale 1ns/1ps

// Integration step 2: CSR + CE + FIFOs + FSM with simple device
// Uses the internal simplified qspi_device to supply 0xFF data.
module int_csr_ce_fsm_tb;
  reg clk; reg resetn;

  // APB
  reg        psel; reg penable; reg pwrite; reg [11:0] paddr; reg [31:0] pwdata; reg [3:0] pstrb;
  wire [31:0] prdata; wire pready; wire pslverr;

  // QSPI pads
  wire sclk; wire cs_n; wire [3:0] io;

  // CSR <-> CE wires
  wire enable_w, xip_en_w, quad_en_w, cpol_w, cpha_w, cmd_start_w, dma_en_w, mode_en_w;
  wire [2:0] clk_div_w; wire cs_auto_w;
  wire [1:0] cmd_lanes_w, addr_lanes_w, data_lanes_w, addr_bytes_w; wire [3:0] dummy_cycles_w;
  wire is_write_w; wire [7:0] opcode_w, mode_bits_w; wire [31:0] cmd_addr_w, cmd_len_w; wire [7:0] extra_dummy_w;
  wire cmd_trigger_clr_w;

  // FIFOs
  wire [31:0] fifo_tx_data_csr_w; wire fifo_tx_we_csr_w; wire [31:0] fifo_tx_rd_data_w; wire fifo_tx_rd_en_w;
  wire fifo_tx_full_w, fifo_tx_empty_w; wire [4:0] fifo_tx_level_w;
  wire fifo_rx_re_csr_w; wire [31:0] fifo_rx_rd_data_w; wire fifo_rx_full_w, fifo_rx_empty_w; wire [4:0] fifo_rx_level_w;

  // CE <-> FSM
  wire fsm_start_w, fsm_done_w;
  wire [31:0] fsm_rx_data_w; wire fsm_rx_wen_w; wire fsm_tx_ren_w;

  // CSR
  csr u_csr (
    .pclk(clk), .presetn(resetn),
    .psel(psel), .penable(penable), .pwrite(pwrite), .paddr(paddr), .pwdata(pwdata), .pstrb(pstrb),
    .prdata(prdata), .pready(pready), .pslverr(pslverr),
    .enable_o(enable_w), .xip_en_o(xip_en_w), .quad_en_o(quad_en_w), .cpol_o(cpol_w), .cpha_o(cpha_w), .lsb_first_o(),
    .cmd_start_o(cmd_start_w), .dma_en_o(dma_en_w), .mode_en_o(mode_en_w), .hold_en_o(), .wp_en_o(),
    .cmd_trigger_clr_i(cmd_trigger_clr_w),
    .clk_div_o(clk_div_w), .cs_auto_o(cs_auto_w), .cs_level_o(), .cs_delay_o(),
    .xip_addr_bytes_o(), .xip_data_lanes_o(), .xip_dummy_cycles_o(), .xip_cont_read_o(), .xip_mode_en_o(), .xip_write_en_o(),
    .xip_read_op_o(), .xip_mode_bits_o(), .xip_write_op_o(),
    .cmd_lanes_o(cmd_lanes_w), .addr_lanes_o(addr_lanes_w), .data_lanes_o(data_lanes_w), .addr_bytes_o(addr_bytes_w),
    .mode_en_cfg_o(), .dummy_cycles_o(dummy_cycles_w), .is_write_o(is_write_w), .opcode_o(opcode_w), .mode_bits_o(mode_bits_w),
    .cmd_addr_o(cmd_addr_w), .cmd_len_o(cmd_len_w), .extra_dummy_o(extra_dummy_w),
    .burst_size_o(), .dma_dir_o(), .incr_addr_o(), .dma_addr_o(), .dma_len_o(),
    .fifo_tx_data_o(fifo_tx_data_csr_w), .fifo_tx_we_o(fifo_tx_we_csr_w),
    .fifo_rx_data_i(fifo_rx_rd_data_w), .fifo_rx_re_o(fifo_rx_re_csr_w),
    .int_en_o(),
    .cmd_done_set_i(fsm_done_w), .dma_done_set_i(1'b0), .err_set_i(1'b0), .fifo_tx_empty_set_i(1'b0), .fifo_rx_full_set_i(1'b0),
    .busy_i(1'b0), .xip_active_i(1'b0), .cmd_done_i(1'b0), .dma_done_i(1'b0),
    .tx_level_i(fifo_tx_level_w[3:0]), .rx_level_i(fifo_rx_level_w[3:0]), .tx_empty_i(fifo_tx_empty_w), .rx_full_i(fifo_rx_full_w),
    .timeout_i(1'b0), .overrun_i(1'b0), .underrun_i(1'b0), .axi_err_i(1'b0), .irq()
  );

  // CE
  cmd_engine #(.ADDR_WIDTH(32)) u_ce (
    .clk(clk), .resetn(resetn), .cmd_start_i(cmd_start_w), .cmd_trigger_clr_o(cmd_trigger_clr_w), .cmd_done_set_o(), .busy_o(),
    .cmd_lanes_i(cmd_lanes_w), .addr_lanes_i(addr_lanes_w), .data_lanes_i(data_lanes_w), .addr_bytes_i(addr_bytes_w),
    .mode_en_i(mode_en_w), .dummy_cycles_i(dummy_cycles_w), .extra_dummy_i(extra_dummy_w), .is_write_i(is_write_w),
    .opcode_i(opcode_w), .mode_bits_i(mode_bits_w), .cmd_addr_i(cmd_addr_w), .cmd_len_i(cmd_len_w),
    .quad_en_i(quad_en_w), .cs_auto_i(cs_auto_w), .xip_cont_read_i(1'b0), .clk_div_i(clk_div_w), .cpol_i(cpol_w), .cpha_i(cpha_w),
    .start_o(fsm_start_w), .done_i(fsm_done_w),
    .cmd_lanes_o(), .addr_lanes_o(), .data_lanes_o(), .addr_bytes_o(), .mode_en_o(), .dummy_cycles_o(), .dir_o(),
    .quad_en_o(), .cs_auto_o(), .xip_cont_read_o(), .opcode_o(), .mode_bits_o(), .addr_o(), .len_o(), .clk_div_o(), .cpol_o(), .cpha_o()
  );

  // FIFOs
  fifo_tx #(.WIDTH(32), .DEPTH(16)) u_ftx (
    .clk(clk), .resetn(resetn),
    .wr_en_i(fifo_tx_we_csr_w), .wr_data_i(fifo_tx_data_csr_w),
    .rd_en_i(fifo_tx_rd_en_w), .rd_data_o(fifo_tx_rd_data_w),
    .full_o(fifo_tx_full_w), .empty_o(fifo_tx_empty_w), .level_o(fifo_tx_level_w)
  );
  fifo_rx #(.WIDTH(32), .DEPTH(16)) u_frx (
    .clk(clk), .resetn(resetn),
    .wr_en_i(fsm_rx_wen_w), .wr_data_i(fsm_rx_data_w),
    .rd_en_i(fifo_rx_re_csr_w), .rd_data_o(fifo_rx_rd_data_w),
    .full_o(fifo_rx_full_w), .empty_o(fifo_rx_empty_w), .level_o(fifo_rx_level_w)
  );

  // FSM
  qspi_fsm u_fsm (
    .clk(clk), .resetn(resetn), .start(fsm_start_w), .done(fsm_done_w),
    .cmd_lanes_sel(cmd_lanes_w), .addr_lanes_sel(addr_lanes_w), .data_lanes_sel(data_lanes_w), .addr_bytes_sel(addr_bytes_w),
    .mode_en(1'b0), .dummy_cycles(dummy_cycles_w), .dir(1'b1), .quad_en(1'b0), .cs_auto(1'b1), .cs_delay(2'b00), .xip_cont_read(1'b0),
    .cmd_opcode(opcode_w), .mode_bits(8'h00), .addr(cmd_addr_w), .len_bytes(cmd_len_w),
    .clk_div({29'd0, clk_div_w}), .cpol(cpol_w), .cpha(cpha_w),
    .tx_data_fifo(fifo_tx_rd_data_w), .tx_empty(fifo_tx_empty_w), .tx_ren(fifo_tx_rd_en_w),
    .rx_data_fifo(fsm_rx_data_w), .rx_wen(fsm_rx_wen_w), .rx_full(fifo_rx_full_w),
    .sclk(sclk), .cs_n(cs_n), .io0(io[0]), .io1(io[1]), .io2(io[2]), .io3(io[3])
  );

  // Simple device
  qspi_device dev (
    .qspi_sclk(sclk), .qspi_cs_n(cs_n), .qspi_io0(io[0]), .qspi_io1(io[1]), .qspi_io2(io[2]), .qspi_io3(io[3])
  );

  // Clock/reset
  initial clk=0; always #5 clk=~clk; initial resetn=0;

  // Debug capture
  reg seen_word; reg [31:0] last_data;
  always @(posedge clk) begin
    if (!resetn) begin seen_word<=1'b0; last_data<=32'h0; end
    else if (fsm_rx_wen_w) begin
      last_data <= fsm_rx_data_w;
      seen_word <= 1'b1;
      $display("[int2] rx_wen data=%08h time=%0t", fsm_rx_data_w, $time);
    end
  end
  integer sclk_edges;
  reg cs_n_q;
  always @(posedge clk) begin
    cs_n_q <= cs_n;
    if (!cs_n && (sclk===1'b0 || sclk===1'b1)) begin
      // crude edge detect by comparing sampled sclk to previous sample
    end
  end

  // APB helpers
  task apb_write(input [11:0] addr, input [31:0] data);
  begin @(posedge clk); psel<=1;penable<=0;pwrite<=1;paddr<=addr;pwdata<=data;pstrb<=4'hF; @(posedge clk); penable<=1; @(posedge clk);
        psel<=0;penable<=0;pwrite<=0;paddr<=0;pwdata<=0;pstrb<=0; end endtask
  task apb_read(input [11:0] addr, output [31:0] data);
  begin @(posedge clk); psel<=1;penable<=0;pwrite<=0;paddr<=addr; @(posedge clk); penable<=1; @(posedge clk); data=prdata; psel<=0; penable<=0; paddr<=0; end endtask

  // CSR addrs
  localparam CTRL=12'h004, CLKDIV=12'h014, CS_CTRL=12'h018, CMD_CFG=12'h024, CMD_OP=12'h028, CMD_ADDR=12'h02C, CMD_LEN=12'h030, FIFO_RX=12'h048, FIFO_STAT=12'h04C;

  integer i; reg [31:0] d;
  initial begin
    psel=0;penable=0;pwrite=0;paddr=0;pwdata=0;pstrb=0; repeat(10) @(posedge clk); resetn=1;
    // Mode0, slow clock, CS auto
    apb_write(CTRL,   32'h0000_0001);
    apb_write(CLKDIV, 32'h0000_0004);
    apb_write(CS_CTRL,32'h0000_0001);
    // 0x03 read 4B @ 0
    apb_write(CMD_CFG,32'h0000_0040);
    apb_write(CMD_OP, 32'h0000_0003);
    apb_write(CMD_ADDR,32'h0000_0000);
    apb_write(CMD_LEN, 32'h0000_0004);
    apb_write(CTRL,   32'h0000_0101);
    // wait capture event
    for (i=0;i<20000 && !seen_word;i=i+1) @(posedge clk);
    if (!seen_word) $fatal(1, "int_csr_ce_fsm: no RX word observed");
    if (last_data !== 32'h7FFF_FFFF && last_data !== 32'hFFFF_FFFF)
      $fatal(1, "int_csr_ce_fsm: expected 7FFFFFFF/FFFFFFFF got %h", last_data);
    $display("CSR+CE+FSM integration test passed");
    $finish;
  end

  // Global timeout to prevent stalls
  initial begin
    #1_000_000; // 1 ms cutoff
    $display("[int_csr_ce_fsm_tb] Global timeout reached — finishing.");
    $finish;
  end
endmodule
